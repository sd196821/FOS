`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:09:36 10/07/2015 
// Design Name: 
// Module Name:    SC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "BRAN.cfg"
`define REG_WIDTH 7
module SC(
			input [`REG_WIDTH-1:0] srs1,
			input [`REG_WIDTH-1:0] srs2,
			input [`REG_WIDTH-1:0] srs3,
			input [`REG_WIDTH-1:0] srd,
			
			input [X_LEN-1:0]rd_data,
			output 
			
			input clk,
			input 
			);


endmodule
