`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:32:38 10/02/2015 
// Design Name: 
// Module Name:    FETCH 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "BEAN.cfg"
module FETCH(
				input reg [`XPR_LEN-1:0] pc,
				output reg [`XPR_LEN-1:0] command,
				input clk
				);

//always @(posedge clk)
//begin

//end

endmodule
